interface dff_intf (input logic clk);
  logic reset;
  logic d;
  logic q;
endinterface
